LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY memory IS
	PORT (
		dir : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
		data : OUT STD_LOGIC_VECTOR (93 DOWNTO 0));
END memory;

ARCHITECTURE Behavioral OF memory IS

BEGIN
	PROCESS (dir)
	BEGIN
		-- DATA FORMAT
		-- |    PRUEBA    |VF| Ins |                LIGA                 |
		--  P4 P3 P2 P1 P0 VF I1 I0 L11 L10 L9 L8 L7 L6 L5 L4 L3 L2 L1 L0 nCRI EB1 EB0 nWB EA1 EA0 nWA selbus UPA9 UPA8 UPA7 UPA6 UPA5 UPA4 UPA3 UPA2 UPA1 UPA0 nOEUPA nDUPA selmux nEX2 nEX1 nEX0 X2 X1 X0 EnaY nERA2 nERA1 nERA0 RA2 RA1 RA0 nEAP2 nEAP1 nEAP0 AP2 AP1 AP0 nEPC2 nEPC1 nEPC0 PC2 PC1 PC0 nCBD nAS nRW BD DINT HINT SET_IRQ SET_XIRQ B9 B8 B7 B6 B5 B4 B3 B2 B1 B0 CC CN CV CZ CI CH CX CS nHB ACCSEC

		-- Cadena por default: "00000" & "0" & "00" & "000000000000" & "10010010000000000011011100001110001110001110001110000000000000000000000010"

		--if(dir=    X"000") then data <= "00000" & "0" & "00" & "000000000000" & "10010010000000000011011100001110001110001110001110000000000000000000000010";
		--elsif(dir= X"001") then data <= "00000" & "0" & "00" & "000000000000" & "00000000000000000000000000000000000000000000000000000000000000000000000000"; 
		IF (dir = X"008") THEN
			data <= "0000000000000000000010010010000000000011011100001110001110000110000110000000000000000000000010";
		ELSIF (dir = X"009") THEN
			data <= "0000000000000000000000010010000000000011011100001110001110001110011010000000000000000000000010";
		ELSIF (dir = X"00A") THEN
			data <= "0000001000000000000010010010000000000011011100001110001110001110001110000000000000000000000010";
			--instrucciones
		ELSIF (dir = X"860") THEN
			data <= "0000000000000000000010010010000000000011011100001110001110000110000110000000000000000000000010";
		ELSIF (dir = X"861") THEN
			data <= "0000000000000000000010010100000000000011011100001110001110001110011010000000000000000000000010";
		ELSIF (dir = X"862") THEN
			data <= "0111111100000000000010010010000000000011011100001110001110001110001110000000010011000111000010";
		ELSIF (dir = X"863") THEN
			data <= "1100000100000000100110010010000000000011011100001110001110000110000110000000000000000000000010";
		ELSIF (dir = X"C60") THEN
			data <= "0000000000000000000010010010000000000011011100001110001110000110000110000000000000000000000010";
		ELSIF (dir = X"C61") THEN
			data <= "0000000000000000000010010100000000000011011100001110001110001110011010000000000000000000000010";
		ELSIF (dir = X"C62") THEN
			data <= "0111111100000000000010010010000000000011011100001110001110001110001110000000100101000111000010";
		ELSIF (dir = X"C63") THEN
			data <= "1100000100000000100110010010000000000011011100001110001110000110000110000000000000000000000010";
		ELSIF (dir = X"CE0") THEN
			data <= "0000000000000000000010010010000000000011011100001110001110000110000110000000000000000000000010";
		ELSIF (dir = X"CE1") THEN
			data <= "0000000000000000000010010010000000000011011001101110001110001110011010000000000000000000000010";
		ELSIF (dir = X"CE2") THEN
			data <= "0111111100000000000010010010000000000011011100001110001110001110001110000000110111000111000010";
		ELSIF (dir = X"CE3") THEN
			data <= "1100000100000000100110010010000000000011011100001110001110000110000110000000000000000000000010";
		ELSIF (dir = X"A50") THEN
			data <= "0000000000000000000010010010000000000011001100001110001110001110000110000000000000000000000010";
		ELSIF (dir = X"A51") THEN
			data <= "0000000000000000000010010010000000000011011100001100111110001110001010000000000000000000000010";
		ELSIF (dir = X"A52") THEN
			data <= "0111111100000000000010010010000000000011011100001100001110001110001110000000000000011000000010";
		ELSIF (dir = X"A53") THEN
			data <= "1100000100000000100110010010000000000011011100001110001110000110000110000000000000000000000010";
		ELSIF (dir = X"200") THEN
			data <= "0000000000000000000010010010000000000011011100001100111110000110000110000000000000000000000000";
		ELSIF (dir = X"201") THEN
			data <= "0000000000000000000010010010000011011111011100001110001110001110011010000000000000000000000010";
		ELSIF (dir = X"202") THEN
			data <= "0000000000000000000010010010001000011011111100001110001110001100001110000000000000000000000010";
		ELSIF (dir = X"203") THEN
			data <= "0000010100100000100010010010000000000000011100001110001110001100111110000000000000001000000010";
		ELSIF (dir = X"204") THEN
			data <= "0000000000000000000010010011001000011111011100001110001110001010001110000000000000000000000010";
		ELSIF (dir = X"205") THEN
			data <= "0000000000000000000010010010000000000000011100001110001110001011001110000000000000000000000010";
		ELSIF (dir = X"206") THEN
			data <= "0000000000000000000010010010000000000011011100001100001110001110001110000000000000011000000000";
		ELSIF (dir = X"207") THEN
			data <= "0111111100000000000010010010000000000011011100001110001110000110000110000000000000000000000010";
		ELSIF (dir = X"208") THEN
			data <= "0100000100000000100110010011001010011111011100001110001110001010001110000000000000000000000010";
		ELSIF (dir = X"260") THEN
			data <= "1001000100100000000110010010000000000011011100001100111110000110000110000000000000000000000000";
		ELSIF (dir = X"261") THEN
			data <= "0111111100000000000010010010000000000011011100001110001110001110011110000000000000000000000010";
		ELSIF (dir = X"262") THEN
			data <= "1100000100000000100110010010000000000011011100001110001110000110000110000000000000000000000010";
		ELSIF (dir = X"270") THEN
			data <= "1001010100100000000110010010000000000011011100001100111110000110000110000000000000000000000000";
		ELSIF (dir = X"271") THEN
			data <= "0111111100000000000010010010000000000011011100001110001110001110011110000000000000000000000010";
		ELSIF (dir = X"272") THEN
			data <= "1100000100000000100110010010000000000011011100001110001110000110000110000000000000000000000010";
		ELSIF (dir = X"240") THEN
			data <= "1000000100100000000110010010000000000011011100001100111110000110000110000000000000000000000000";
		ELSIF (dir = X"241") THEN
			data <= "0111111100000000000010010010000000000011011100001110001110001110011110000000000000000000000010";
		ELSIF (dir = X"242") THEN
			data <= "1100000100000000100110010010000000000011011100001110001110000110000110000000000000000000000010";
		ELSIF (dir = X"250") THEN
			data <= "1000010100100000000110010010000000000011011100001100111110000110000110000000000000000000000000";
		ELSIF (dir = X"251") THEN
			data <= "0111111100000000000010010010000000000011011100001110001110001110011110000000000000000000000010";
		ELSIF (dir = X"252") THEN
			data <= "1100000100000000100110010010000000000011011100001110001110000110000110000000000000000000000010";
		ELSIF (dir = X"2B0") THEN
			data <= "1001110100100000000110010010000000000011011100001100111110000110000110000000000000000000000000";
		ELSIF (dir = X"2B1") THEN
			data <= "0111111100000000000010010010000000000011011100001110001110001110011110000000000000000000000010";
		ELSIF (dir = X"2B2") THEN
			data <= "1100000100000000100110010010000000000011011100001110001110000110000110000000000000000000000010";
		ELSIF (dir = X"2A0") THEN
			data <= "1001100100100000000110010010000000000011011100001100111110000110000110000000000000000000000000";
		ELSIF (dir = X"2A1") THEN
			data <= "0111111100000000000010010010000000000011011100001110001110001110011110000000000000000000000010";
		ELSIF (dir = X"2A2") THEN
			data <= "1100000100000000100110010010000000000011011100001110001110000110000110000000000000000000000010";
		ELSIF (dir = X"db0") THEN
			data <= "0000000000000000000010010010000000000011011100001110001110000110000110000000000000000000000010";
		ELSIF (dir = X"db1") THEN
			data <= "0000000000000000000010010010000000000011011100001100111110001110011010000000000000000000000010";
		ELSIF (dir = X"db2") THEN
			data <= "0000000000000000000010010010000000000011011100000110001110001110000110000000000000000000000010";
		ELSIF (dir = X"db3") THEN
			data <= "0000000000000000000010011110001000010111111100001110001110001110001010000000000000000000000011";
		ELSIF (dir = X"db4") THEN
			data <= "0111111100000000000010010100000000000000011100001110001110001110001110000000000000001111000010";
		ELSIF (dir = X"db5") THEN
			data <= "1100000100000000100110010010000000000011011100001110001110000110000110000000000000000000000010";
		ELSIF (dir = X"8C0") THEN
			data <= "0000000000000000000010010010000000000011011100001110001110000110000110000000000000000000000010";
		ELSIF (dir = X"8C1") THEN
			data <= "0000000000000000000010010010000000000011011100001100111110001110011010000000000000000000000010";
		ELSIF (dir = X"8C2") THEN
			data <= "0000000000000000000010010010000011011111011100001100001110001110001110000000000000000000000010";
		ELSIF (dir = X"8C3") THEN
			data <= "0000000000000000000010010010000001011011111000001110001110001110001110000000000000001111000010";
		ELSIF (dir = X"8C3") THEN
			data <= "0111111100000000000010010010000001011011111000001110001110001110001110000000000000001111000010";
		ELSIF (dir = X"8C4") THEN
			data <= "1100000100000000100110010010000000000011011100001110001110000110000110000000000000000000000010";
		ELSIF (dir = X"080") THEN
			data <= "0000000000000000000010010010000000000011011100101110001110001110001110000000000000000000000010";
		ELSIF (dir = X"081") THEN
			data <= "0111111100000000000010010010000000000011011100001110001110001110001110000000000110000001000010";
		ELSIF (dir = X"082") THEN
			data <= "1100000100000000100110010010000000000011011100001110001110000110000110000000000000000000000010";
		ELSIF (dir = X"AD0") THEN
			data <= "0000000000100000000111111110001000000111111100001110001110001110001110000000000000000000000010";
		ELSIF (dir = X"AD1") THEN
			data <= "0111111100000000000010010010000000000000011001101110001110001110001110000000000000001111000010";
		ELSIF (dir = X"AD2") THEN
			data <= "1100000100000000100110010010000000000011011100001110001110000110000110000000000000000000000010";
		ELSIF (dir = X"7E0") THEN
			data <= "0000000000000000000010010010000000000011011100001110001110000110000110000000000000000000000010";
		ELSIF (dir = X"7E1") THEN
			data <= "0000000000000000000010010010000000000011011100001011001110001110011011000000000000000000000010";
		ELSIF (dir = X"7E2") THEN
			data <= "0000000000000000000010010010000000000011011100001110001110000110000110000000000000000000000010";
		ELSIF (dir = X"7E3") THEN
			data <= "0000000000000000000010010010000000000011011100001100111110001110001010000000000000000000000010";
		ELSIF (dir = X"7E4") THEN
			data <= "0000000000000000000010010010000000000011011100001000001110001001011110000000000000000000000010";
		ELSIF (dir = X"7E5") THEN
			data <= "0111111100000000000010010010000000000011011100001110001110001110001110000000000000000000000010";
		ELSIF (dir = X"7E6") THEN
			data <= "1100000100000000100110010010000000000011011100001110001110000110000110000000000000000000000010";
		ELSIF (dir = X"e00") THEN
			data <= "0000000000000000000010010010000000000011011100001110001110000110000110000000000000000000000010";
		ELSIF (dir = X"e01") THEN
			data <= "0000000000000000000010010010000011011111011100001110001110001110011010000000000000000000000010";
		ELSIF (dir = X"e02") THEN
			data <= "0000000000000000000010010010001000011011111100001110001110001110001110000000000000000000000010";
		ELSIF (dir = X"e03") THEN
			data <= "0000000000000000000010010010000000000000011100001100111110001110001110000000000000001000000010";
		ELSIF (dir = X"e04") THEN
			data <= "0000000000000000000010010011000000011111011100001010001110001110001110000000000000000000000010";
		ELSIF (dir = X"e05") THEN
			data <= "0000000000000000000010010010000000000000011100001011001110001110001110000000000000000000000010";
		ELSIF (dir = X"e06") THEN
			data <= "0000000000000000000010010010000000000011011100000110001110001110000110000000000000000000000010";
		ELSIF (dir = X"e07") THEN
			data <= "0000000000000000000011110010000001100011111100001110001110001110001010000000000000000000000010";
		ELSIF (dir = X"e08") THEN
			data <= "0111111100000000000010100010000000000000011100001110001110001110001110000000000000001111010010";
		ELSIF (dir = X"e09") THEN
			data <= "1100000100000000100110010010000000000011011100001110001110000110000110000000000000000000000010";
		ELSIF (dir = X"ab0") THEN
			data <= "0000000000000000000010010010000000000011011100001110001110000110000110000000000000000000000010";
		ELSIF (dir = X"ab1") THEN
			data <= "0000000000000000000010010010000011011111011100001110001110001110011010000000000000000000000010";
		ELSIF (dir = X"ab2") THEN
			data <= "0000000000000000000010010010000000011011111000001110001110001110001110000000000000000000000010";
		ELSIF (dir = X"ab3") THEN
			data <= "0000000000000000000010010010000000000000011100001100111110001110001110000000000000001000000010";
		ELSIF (dir = X"ab4") THEN
			data <= "0000000000000000000010010011000000001011011100001010001110001110001110000000000000000000000010";
		ELSIF (dir = X"ab5") THEN
			data <= "0000000000000000000010010010000000000000011100001011001110001110001110000000000000000000000010";
		ELSIF (dir = X"ab6") THEN
			data <= "0000000000000000000010010010000000000011011100000110001110001110000110000000000000000000000010";
		ELSIF (dir = X"ab7") THEN
			data <= "0000000000000000000010011110000000010111111100001110001110001110001010000000000000000000000010";
		ELSIF (dir = X"ab8") THEN
			data <= "0111111100000000000010010100000000000000011100001110001110001110001110000000000000001111010010";
		ELSIF (dir = X"ab9") THEN
			data <= "1100000100000000100110010010000000000011011100001110001110000110000110000000000000000000000010";
		ELSE
			data <= "0000000000000000100010010010000000000011011100001110001110001110001110000000000000000000000010"; -- Default
		END IF;
	END PROCESS;
END Behavioral;